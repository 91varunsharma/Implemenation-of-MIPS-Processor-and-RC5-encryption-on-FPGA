----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:12:06 12/05/2016 
-- Design Name: 
-- Module Name:    IFetch - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

Entity IFetch is
    Port (
           NextPC      : in  STD_LOGIC_VECTOR (31 downto 0);
           --PC          : out  STD_LOGIC_VECTOR (31 downto 0);
           Instruction : out  STD_LOGIC_VECTOR (31 downto 0));
End IFetch;


architecture Behavioral of IFetch is
    
--SIGNAL Program_Counter : STD_LOGIC_VECTOR (31 downto 0);
-- change array index to 1023 later
Type IMemory IS ARRAY (0 to 589) of STD_LOGIC_VECTOR(31 downto 0);

 CONSTANT IMem : IMemory:=IMemory'(X"00006010",X"00006810",X"00000810",X"00001010",X"040e004d",X"040a0019",X"040b0003",X"04140001",
X"04110000",X"04120028",X"00000000",X"00000000",X"00000000",X"1e2f0000",X"00222810",X"00af2810",
X"30000034",X"00060810",X"22210000",X"00224810",X"1e500000",X"02093810",X"0d29001f",X"0007b010",
X"0009c010",X"300000a2",X"00174010",X"00081010",X"22420000",X"294c000a",X"058c0001",X"06310001",
X"296d000d",X"05ad0001",X"06520001",X"280e001d",X"09ce0001",X"3000000d",X"00000000",X"00000000",
X"04110000",X"040c0000",X"30000020",X"00000000",X"00000000",X"00000000",X"04120028",X"040d0000",
X"30000023",X"00000000",X"00000000",X"00000000",X"0415ffff",X"16b5001d",X"00b5a812",X"1ab5001d",
X"14a50003",X"00b53013",X"30000011",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
X"00000000",X"00006810",X"00002010",X"04030019",X"1c010032",X"1c020033",X"040b0000",X"1d6c0000",
X"002c0810",X"056b0001",X"04840001",X"1d6c0000",X"004c1010",X"00000000",X"00000000",X"04140002",
X"0022f013",X"0022f812",X"03df2811",X"0005b010",X"0c4d001f",X"000dc010",X"300000a2",X"00173810",
X"056b0001",X"04840001",X"1d6c0000",X"00ec0810",X"0022f013",X"0022f812",X"03df3011",X"0006b010",
X"0c2d001f",X"000dc010",X"04140004",X"300000a2",X"00174010",X"056b0001",X"04840001",X"1d6c0000",
X"010c1010",X"20010034",X"20020035",X"28640004",X"3000004f",X"00000000",X"00000000",X"00000000",
X"00006810",X"04030002",X"04040019",X"1c010037",X"1c020038",X"040b0019",X"1d6c0000",X"04140003",
X"004c1011",X"0002b010",X"0c2d001f",X"000dc010",X"300000e4",X"00174010",X"0101f013",X"0101f812",
X"03df3011",X"00061010",X"08840001",X"096b0001",X"1d6c0000",X"002c0811",X"0001b010",X"0c4d001f",
X"000dc010",X"04140005",X"300000e4",X"00173810",X"00e2f013",X"00e2f812",X"03df2811",X"00050810",
X"28640004",X"08840001",X"096b0001",X"30000076",X"00000000",X"096b0001",X"1d6c0000",X"004c1011",
X"096b0001",X"1d6c0000",X"002c0811",X"20010039",X"2002003a",X"3000024d",X"00000000",X"00000000",
X"00000000",X"00000000",X"0415ffff",X"00009810",X"2a780197",X"06730001",X"2a780080",X"06730001",
X"2a780087",X"06730001",X"2a78008e",X"06730001",X"2a780095",X"06730001",X"2a78009c",X"06730001",
X"2a7800a3",X"06730001",X"2a7800aa",X"06730001",X"2a7800b1",X"06730001",X"2a7800b8",X"06730001",
X"2a7800bf",X"06730001",X"2a7800c6",X"06730001",X"2a7800cd",X"06730001",X"2a7800d4",X"06730001",
X"2a7800db",X"06730001",X"2a7800e2",X"06730001",X"2a7800e9",X"06730001",X"2a7800f0",X"06730001",
X"2a7800f7",X"06730001",X"2a7800fe",X"06730001",X"2a780105",X"06730001",X"2a78010c",X"06730001",
X"2a780113",X"06730001",X"2a78011a",X"06730001",X"2a780121",X"06730001",X"2a780128",X"06730001",
X"2a78012f",X"06730001",X"2a780136",X"06730001",X"2a78013d",X"06730001",X"2a780144",X"06730001",
X"2a78014b",X"06730001",X"2a780152",X"00000000",X"0415ffff",X"00009810",X"2a780155",X"06730001",
X"2a78014c",X"06730001",X"2a780141",X"06730001",X"2a780136",X"06730001",X"2a78012b",X"06730001",
X"2a780120",X"06730001",X"2a780115",X"06730001",X"2a78010a",X"06730001",X"2a7800ff",X"06730001",
X"2a7800f4",X"06730001",X"2a7800e9",X"06730001",X"2a7800de",X"06730001",X"2a7800d3",X"06730001",
X"2a7800c8",X"06730001",X"2a7800bd",X"06730001",X"2a7800b2",X"06730001",X"2a7800a7",X"06730001",
X"2a78009c",X"06730001",X"2a780091",X"06730001",X"2a780086",X"06730001",X"2a78007b",X"06730001",
X"2a780070",X"06730001",X"2a780065",X"06730001",X"2a78005a",X"06730001",X"2a78004f",X"06730001",
X"2a780044",X"06730001",X"2a780039",X"06730001",X"2a78002e",X"06730001",X"2a780023",X"06730001",
X"2a780018",X"06730001",X"2a78000d",X"06730001",X"2a780002",X"00000000",X"00000000",X"16b5001f",
X"02d5a812",X"1ab5001f",X"16d60001",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",
X"16b5001e",X"02d5a812",X"1ab5001e",X"16d60002",X"02d5b813",X"30000242",X"00000000",X"00000000",
X"00000000",X"16b5001d",X"02d5a812",X"1ab5001d",X"16d60003",X"02d5b813",X"30000242",X"00000000",
X"00000000",X"00000000",X"16b5001c",X"02d5a812",X"1ab5001c",X"16d60004",X"02d5b813",X"30000242",
X"00000000",X"00000000",X"00000000",X"16b5001b",X"02d5a812",X"1ab5001b",X"16d60005",X"02d5b813",
X"30000242",X"00000000",X"00000000",X"00000000",X"16b5001a",X"02d5a812",X"1ab5001a",X"16d60006",
X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50019",X"02d5a812",X"1ab50019",
X"16d60007",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50018",X"02d5a812",
X"1ab50018",X"16d60008",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50017",
X"02d5a812",X"1ab50017",X"16d60009",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",
X"16b50016",X"02d5a812",X"1ab50016",X"16d6000a",X"02d5b813",X"30000242",X"00000000",X"00000000",
X"00000000",X"16b50015",X"02d5a812",X"1ab50015",X"16d6000b",X"02d5b813",X"30000242",X"00000000",
X"00000000",X"00000000",X"16b50014",X"02d5a812",X"1ab50014",X"16d6000c",X"02d5b813",X"30000242",
X"00000000",X"00000000",X"00000000",X"16b50013",X"02d5a812",X"1ab50013",X"16d6000d",X"02d5b813",
X"30000242",X"00000000",X"00000000",X"00000000",X"16b50012",X"02d5a812",X"1ab50012",X"16d6000e",
X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50011",X"02d5a812",X"1ab50011",
X"16d6000f",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50010",X"02d5a812",
X"1ab50010",X"16d60010",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b5000f",
X"02d5a812",X"1ab5000f",X"16d60011",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",
X"16b5000e",X"02d5a812",X"1ab5000e",X"16d60012",X"02d5b813",X"30000242",X"00000000",X"00000000",
X"00000000",X"16b5000d",X"02d5a812",X"1ab5000d",X"16d60013",X"02d5b813",X"30000242",X"00000000",
X"00000000",X"00000000",X"16b5000c",X"02d5a812",X"1ab5000c",X"16d60014",X"02d5b813",X"30000242",
X"00000000",X"00000000",X"00000000",X"16b5000b",X"02d5a812",X"1ab5000b",X"16d60015",X"02d5b813",
X"30000242",X"00000000",X"00000000",X"00000000",X"16b5000a",X"02d5a812",X"1ab5000a",X"16d60016",
X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50009",X"02d5a812",X"1ab50009",
X"16d60017",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50008",X"02d5a812",
X"1ab50008",X"16d60018",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50007",
X"02d5a812",X"1ab50007",X"16d60019",X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",
X"16b50006",X"02d5a812",X"1ab50006",X"16d6001a",X"02d5b813",X"30000242",X"00000000",X"00000000",
X"00000000",X"16b50005",X"02d5a812",X"1ab50005",X"16d6001b",X"02d5b813",X"30000242",X"00000000",
X"00000000",X"00000000",X"16b50004",X"02d5a812",X"1ab50004",X"16d6001c",X"02d5b813",X"30000242",
X"00000000",X"00000000",X"00000000",X"16b50003",X"02d5a812",X"1ab50003",X"16d6001d",X"02d5b813",
X"30000242",X"00000000",X"00000000",X"00000000",X"16b50002",X"02d5a812",X"1ab50002",X"16d6001e",
X"02d5b813",X"30000242",X"00000000",X"00000000",X"00000000",X"16b50001",X"02d5a812",X"1ab50001",
X"16d6001f",X"02d5b813",X"30000242",X"00000000",X"0016b810",X"30000242",X"00000000",X"00000000",
X"00000000",X"00000000",X"04190002",X"2699fdd6",X"07390001",X"2699fe11",X"07390001",X"2699fe35",
X"07390001",X"2699fe1a",X"07390001",X"2699fe3f",X"00000000",X"fc000000");          
     
begin
   
   Instruction <= IMem(conv_integer(NextPC));
   --PC <= NextPC;

End Behavioral;

